`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:22:23 08/25/2014 
// Design Name: 
// Module Name:    lab3dpath 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module lab3dpath(x1,x2,x3,y);
input [9:0] x1,x2,x3;
output [9:0] y;

//complete this module

endmodule
