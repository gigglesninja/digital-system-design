`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:10:52 08/30/2014 
// Design Name: 
// Module Name:    lab4dpath 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module lab4dpath(x1,x2,x3,y,clk);
input clk;
input [9:0] x1,x2,x3;
output [9:0] y;

 
 
endmodule

